module ctrlUnit(
  input wire[6:0] opCode,
  output reg wr_en,m_wr_en, //??????
  output reg[2:0] alu_op  //??????
);

  always @* begin
    if(opCode == 7'b0000001) begin //?????0000001
      wr_en = 1;
      alu_op = 3'b001;  //??????
      m_wr_en = 0;  //??????
    end
    else if(opCode == 7'b0000010) begin //?????? ?????0000010
      wr_en = 0;
      alu_op = 3'b010;  //??????
      m_wr_en = 1;
    end
    else begin
      wr_en = 0;
      alu_op = 3'b000;  //??????
      m_wr_en = 0;  //??????
    end
  
  end
endmodule 
